module tb_uart_tx;
reg clk, rst;
reg tx_start